module cc_saida_ck3hz(
input ea0,
input ea1,
output out
);
buf(out,ea1);
endmodule
